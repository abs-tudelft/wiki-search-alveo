-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

library work;
use work.Axi_pkg.all;
use work.UtilInt_pkg.all;
use work.UtilConv_pkg.all;
use work.UtilMisc_pkg.all;
use work.Array_pkg.all;
use work.vhsnunzip_pkg.all;
use work.vhdmmio_pkg.all;
use work.WordMatch_MMIO_pkg.all;

-------------------------------------------------------------------------------
-- AXI4 compatible top level for Fletcher generated accelerators.
-------------------------------------------------------------------------------
-- Requires an AXI4 port to host memory.
-- Requires an AXI4-lite port from host for MMIO.
-------------------------------------------------------------------------------
-- NOTE: this file is NOT generated by Fletchgen; it has undergone heavy manual
-- optimization to improve performance.
entity WordMatch_AxiTop is
  generic (
    BUS_ADDR_WIDTH              : natural := 64;
    BUS_DATA_WIDTH              : natural := 64;
    BUS_LEN_WIDTH               : natural := 8;
    BUS_READ_INNER_DATA_WIDTH   : natural := 64;
    BUS_READ_BURST_MAX_LEN      : natural := 128;
    BUS_READ_BURST_STEP_LEN     : natural := 8;
    BUS_WRITE_INNER_DATA_WIDTH  : natural := 32;
    BUS_WRITE_BURST_MAX_LEN     : natural := 16;
    BUS_WRITE_BURST_STEP_LEN    : natural := 4
  );
  port (

    -- Bus clock domain.
    bus_clk                     : in  std_logic;
    bus_reset                   : in  std_logic;

    -- Internal clock domain for the decompression and matchers.
    dec_clk                     : in  std_logic;
    dec_reset                   : in  std_logic;

    ---------------------------------------------------------------------------
    -- AXI4 master as Host Memory Interface
    ---------------------------------------------------------------------------
    -- Read address channel
    m_axi_araddr                : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    m_axi_arlen                 : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    m_axi_arvalid               : out std_logic := '0';
    m_axi_arready               : in  std_logic;
    m_axi_arsize                : out std_logic_vector(2 downto 0);

    -- Read data channel
    m_axi_rdata                 : in  std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    m_axi_rresp                 : in  std_logic_vector(1 downto 0);
    m_axi_rlast                 : in  std_logic;
    m_axi_rvalid                : in  std_logic;
    m_axi_rready                : out std_logic := '0';

    -- Write address channel
    m_axi_awvalid               : out std_logic := '0';
    m_axi_awready               : in  std_logic;
    m_axi_awaddr                : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    m_axi_awlen                 : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    m_axi_awsize                : out std_logic_vector(2 downto 0);

    -- Write data channel
    m_axi_wvalid                : out std_logic := '0';
    m_axi_wready                : in  std_logic;
    m_axi_wdata                 : out std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    m_axi_wlast                 : out std_logic;
    m_axi_wstrb                 : out std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);

    -- Write response channel
    m_axi_bvalid                : in  std_logic;
    m_axi_bready                : out std_logic;
    m_axi_bresp                 : in  std_logic_vector(1 downto 0);

    ---------------------------------------------------------------------------
    -- AXI4-lite Slave as MMIO interface
    ---------------------------------------------------------------------------
    -- Write adress channel
    s_axi_awvalid               : in std_logic;
    s_axi_awready               : out std_logic;
    s_axi_awaddr                : in std_logic_vector(31 downto 0);

    -- Write data channel
    s_axi_wvalid                : in std_logic;
    s_axi_wready                : out std_logic;
    s_axi_wdata                 : in std_logic_vector(31 downto 0);
    s_axi_wstrb                 : in std_logic_vector(3 downto 0);

    -- Write response channel
    s_axi_bvalid                : out std_logic;
    s_axi_bready                : in std_logic;
    s_axi_bresp                 : out std_logic_vector(1 downto 0);

    -- Read address channel
    s_axi_arvalid               : in std_logic;
    s_axi_arready               : out std_logic;
    s_axi_araddr                : in std_logic_vector(31 downto 0);

    -- Read data channel
    s_axi_rvalid                : out std_logic;
    s_axi_rready                : in std_logic;
    s_axi_rdata                 : out std_logic_vector(31 downto 0);
    s_axi_rresp                 : out std_logic_vector(1 downto 0)

  );
end WordMatch_AxiTop;

architecture Behavorial of WordMatch_AxiTop is

  -- High-level MMIO register interface provided by vhdMMIO.
  signal mmio_cmd               : wordmatch_mmio_g_cmd_o_type;
  signal mmio_cfg               : wordmatch_mmio_g_cfg_o_type;
  signal mmio_filt              : wordmatch_mmio_g_filt_o_type;
  signal mmio_stat              : wordmatch_mmio_g_stat_i_type;
  signal mmio_start             : std_logic;
  signal mmio_starting          : std_logic;
  signal mmio_done              : std_logic;

  -- Bus signals to convert to AXI.
  signal bus_reset_n            : std_logic;
  signal rd_mst_rreq_addr       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal rd_mst_rreq_len        : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal rd_mst_rreq_valid      : std_logic;
  signal rd_mst_rreq_ready      : std_logic;
  signal rd_mst_rdat_data       : std_logic_vector(BUS_READ_INNER_DATA_WIDTH-1 downto 0);
  signal rd_mst_rdat_last       : std_logic;
  signal rd_mst_rdat_valid      : std_logic;
  signal rd_mst_rdat_ready      : std_logic;
  signal wr_mst_wreq_valid      : std_logic;
  signal wr_mst_wreq_ready      : std_logic;
  signal wr_mst_wreq_addr       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal wr_mst_wreq_len        : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal wr_mst_wdat_valid      : std_logic;
  signal wr_mst_wdat_ready      : std_logic;
  signal wr_mst_wdat_data       : std_logic_vector(BUS_WRITE_INNER_DATA_WIDTH-1 downto 0);
  signal wr_mst_wdat_strobe     : std_logic_vector(BUS_WRITE_INNER_DATA_WIDTH/8-1 downto 0);
  signal wr_mst_wdat_last       : std_logic;
  signal m_axi_awvalid_int      : std_logic;
  signal write_busy             : std_logic;

  -- Typedefs for the internal Fletcher busses.
  type fletcher_read_req is record
    rreq_valid                  : std_logic;
    rreq_addr                   : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    rreq_len                    : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    rdat_ready                  : std_logic;
  end record;

  type fletcher_read_rep is record
    rreq_ready                  : std_logic;
    rdat_valid                  : std_logic;
    rdat_data                   : std_logic_vector(BUS_READ_INNER_DATA_WIDTH-1 downto 0);
    rdat_last                   : std_logic;
  end record;

  type fletcher_read_req_array is array (natural range <>) of fletcher_read_req;
  type fletcher_read_rep_array is array (natural range <>) of fletcher_read_rep;

  type fletcher_write_req is record
    wreq_valid                  : std_logic;
    wreq_addr                   : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    wreq_len                    : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    wdat_valid                  : std_logic;
    wdat_data                   : std_logic_vector(BUS_WRITE_INNER_DATA_WIDTH-1 downto 0);
    wdat_strobe                 : std_logic_vector(BUS_WRITE_INNER_DATA_WIDTH/8-1 downto 0);
    wdat_last                   : std_logic;
  end record;

  type fletcher_write_rep is record
    wreq_ready                  : std_logic;
    wdat_ready                  : std_logic;
  end record;

  -- Signal defs for the internal Fletcher busses.
  signal pages_title_bus_req        : fletcher_read_req;
  signal pages_title_bus_rep        : fletcher_read_rep;
  signal pages_text_bus_req         : fletcher_read_req_array(0 to 2);
  signal pages_text_bus_rep         : fletcher_read_rep_array(0 to 2);
  signal result_title_bus_req       : fletcher_write_req;
  signal result_title_bus_rep       : fletcher_write_rep;
  signal result_count_stats_bus_req : fletcher_write_req;
  signal result_count_stats_bus_rep : fletcher_write_rep;

  -- Page text command/unlock streams.
  signal pages_text_cmd_valid       : std_logic_vector(2 downto 0);
  signal pages_text_cmd_ready       : std_logic_vector(2 downto 0);
  signal pages_text_cmd_idx         : std_logic_vector(127 downto 0);
  signal pages_text_cmd_valuesAddr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal pages_text_cmd_offsetAddr  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal pages_text_cmd_ctrl        : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal pages_text_unl_valid       : std_logic_vector(2 downto 0);
  signal pages_text_unl_ready       : std_logic_vector(2 downto 0);

  -- Match count streams for each of the two partitions.
  signal match_count_part_valid     : std_logic_vector(2 downto 0);
  signal match_count_part_ready     : std_logic_vector(2 downto 0);
  signal match_count_part_amount    : std_logic_vector(47 downto 0);

  -- Arbiter'd match count stream.
  signal match_count_arb_valid      : std_logic;
  signal match_count_arb_ready      : std_logic;
  signal match_count_arb_amount     : std_logic_vector(15 downto 0);
  signal match_count_arb_part       : std_logic_vector(1 downto 0);

  -- Match count stream converted to the bus clock domain.
  signal match_count_xclk_valid     : std_logic;
  signal match_count_xclk_ready     : std_logic;
  signal match_count_xclk_amount    : std_logic_vector(15 downto 0);
  signal match_count_xclk_part      : std_logic_vector(1 downto 0);

  -- Match count stream tagged with the corresponding table indices.
  signal match_count_tagged_valid   : std_logic;
  signal match_count_tagged_ready   : std_logic;
  signal match_count_tagged_amount  : std_logic_vector(15 downto 0);
  signal match_count_tagged_index   : std_logic_vector(19 downto 0);
  signal match_count_tagged_last    : std_logic;

  -- Write command stream.
  signal write_cmd_valid            : std_logic;
  signal write_cmd_ready            : std_logic;
  signal write_cmd_titlePass        : std_logic;
  signal write_cmd_titleDummy       : std_logic;
  signal write_cmd_titleTerm        : std_logic;
  signal write_cmd_intEnable        : std_logic;
  signal write_cmd_intData          : std_logic_vector(31 downto 0);
  signal write_cmd_last             : std_logic;

  -- Page title input command/unlock streams.
  signal pages_title_cmd_valid      : std_logic;
  signal pages_title_cmd_ready      : std_logic;
  signal pages_title_cmd_firstIdx   : std_logic_vector(31 downto 0);
  signal pages_title_cmd_lastidx    : std_logic_vector(31 downto 0);
  signal pages_title_cmd_valuesAddr : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal pages_title_cmd_offsetAddr : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal pages_title_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal pages_title_unl_valid      : std_logic;
  signal pages_title_unl_ready      : std_logic;

  -- Page title input data streams.
  signal pages_title_valid          : std_logic;
  signal pages_title_ready          : std_logic;
  signal pages_title_dvalid         : std_logic;
  signal pages_title_last           : std_logic;
  signal pages_title_length         : std_logic_vector(31 downto 0);
  signal pages_title_count          : std_logic_vector(0 downto 0);
  signal pages_title_chars_valid    : std_logic;
  signal pages_title_chars_ready    : std_logic;
  signal pages_title_chars_dvalid   : std_logic;
  signal pages_title_chars_last     : std_logic;
  signal pages_title_chars_data     : std_logic_vector(7 downto 0);
  signal pages_title_chars_count    : std_logic_vector(0 downto 0);

  -- Result title command/unlock streams.
  signal result_title_cmd_valid     : std_logic;
  signal result_title_cmd_ready     : std_logic;
  signal result_title_cmd_firstIdx  : std_logic_vector(31 downto 0);
  signal result_title_cmd_lastIdx   : std_logic_vector(31 downto 0);
  signal result_title_cmd_valuesAddr: std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal result_title_cmd_offsetAddr: std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal result_title_cmd_ctrl      : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal result_title_unl_valid     : std_logic;
  signal result_title_unl_ready     : std_logic;

  -- Result title output data streams.
  signal result_title_valid         : std_logic;
  signal result_title_ready         : std_logic;
  signal result_title_dvalid        : std_logic;
  signal result_title_last          : std_logic;
  signal result_title_length        : std_logic_vector(31 downto 0);
  signal result_title_count         : std_logic_vector(0 downto 0);
  signal result_title_chars_valid   : std_logic;
  signal result_title_chars_ready   : std_logic;
  signal result_title_chars_dvalid  : std_logic;
  signal result_title_chars_last    : std_logic;
  signal result_title_chars_data    : std_logic_vector(7 downto 0);
  signal result_title_chars_count   : std_logic_vector(0 downto 0);

  -- Result match count & stats command/unlock stream.
  signal result_count_stats_cmd_valid     : std_logic;
  signal result_count_stats_cmd_ready     : std_logic;
  signal result_count_stats_cmd_firstIdx  : std_logic_vector(31 downto 0);
  signal result_count_stats_cmd_lastidx   : std_logic_vector(31 downto 0);
  signal result_count_stats_cmd_addr      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal result_count_stats_unl_valid     : std_logic;
  signal result_count_stats_unl_ready     : std_logic;

  -- Result match count & stats output data stream.
  signal result_count_stats_valid   : std_logic;
  signal result_count_stats_ready   : std_logic;
  signal result_count_stats_data    : std_logic_vector(31 downto 0);
  signal result_count_stats_dvalid  : std_logic;
  signal result_count_stats_last    : std_logic;

begin

  -----------------------------------------------------------------------------
  -- vhdMMIO register file
  -----------------------------------------------------------------------------
  mmio_inst: WordMatch_MMIO
    port map (
      clk                       => bus_clk,
      reset                     => bus_reset,

      g_cmd_o                   => mmio_cmd,
      g_cfg_o                   => mmio_cfg,
      g_filt_o                  => mmio_filt,
      g_stat_i                  => mmio_stat,
      s_start                   => mmio_start,
      s_starting                => mmio_starting,
      s_done                    => mmio_done,

      mmio_awvalid              => s_axi_awvalid,
      mmio_awready              => s_axi_awready,
      mmio_awaddr               => s_axi_awaddr,
      mmio_wvalid               => s_axi_wvalid,
      mmio_wready               => s_axi_wready,
      mmio_wdata                => s_axi_wdata,
      mmio_wstrb                => s_axi_wstrb,
      mmio_bvalid               => s_axi_bvalid,
      mmio_bready               => s_axi_bready,
      mmio_bresp                => s_axi_bresp,
      mmio_arvalid              => s_axi_arvalid,
      mmio_arready              => s_axi_arready,
      mmio_araddr               => s_axi_araddr,
      mmio_rvalid               => s_axi_rvalid,
      mmio_rready               => s_axi_rready,
      mmio_rdata                => s_axi_rdata,
      mmio_rresp                => s_axi_rresp
    );

  -----------------------------------------------------------------------------
  -- AXI interface converter blocks
  -----------------------------------------------------------------------------
  -- Generate active low reset for the converters.
  bus_reset_n <= not bus_reset;

  -- Read datapath.
  axi_read_conv_inst: AxiReadConverter
    generic map (
      ADDR_WIDTH                => BUS_ADDR_WIDTH,
      MASTER_DATA_WIDTH         => BUS_DATA_WIDTH,
      MASTER_LEN_WIDTH          => BUS_LEN_WIDTH,
      SLAVE_DATA_WIDTH          => BUS_READ_INNER_DATA_WIDTH,
      SLAVE_LEN_WIDTH           => BUS_LEN_WIDTH,
      SLAVE_MAX_BURST           => BUS_READ_BURST_MAX_LEN,
      ENABLE_FIFO               => false,
      SLV_REQ_SLICE_DEPTH       => 0,
      SLV_DAT_SLICE_DEPTH       => 0,
      MST_REQ_SLICE_DEPTH       => 0,
      MST_DAT_SLICE_DEPTH       => 0
    )
    port map (
      clk                       => bus_clk,
      reset_n                   => bus_reset_n,
      slv_bus_rreq_addr         => rd_mst_rreq_addr,
      slv_bus_rreq_len          => rd_mst_rreq_len,
      slv_bus_rreq_valid        => rd_mst_rreq_valid,
      slv_bus_rreq_ready        => rd_mst_rreq_ready,
      slv_bus_rdat_data         => rd_mst_rdat_data,
      slv_bus_rdat_last         => rd_mst_rdat_last,
      slv_bus_rdat_valid        => rd_mst_rdat_valid,
      slv_bus_rdat_ready        => rd_mst_rdat_ready,
      m_axi_araddr              => m_axi_araddr,
      m_axi_arlen               => m_axi_arlen,
      m_axi_arvalid             => m_axi_arvalid,
      m_axi_arready             => m_axi_arready,
      m_axi_arsize              => m_axi_arsize,
      m_axi_rdata               => m_axi_rdata,
      m_axi_rlast               => m_axi_rlast,
      m_axi_rvalid              => m_axi_rvalid,
      m_axi_rready              => m_axi_rready
    );

  -- Write datapath.
  axi_write_conv_inst: AxiWriteConverter
    generic map (
      ADDR_WIDTH                => BUS_ADDR_WIDTH,
      MASTER_DATA_WIDTH         => BUS_DATA_WIDTH,
      MASTER_LEN_WIDTH          => BUS_LEN_WIDTH,
      SLAVE_DATA_WIDTH          => BUS_WRITE_INNER_DATA_WIDTH,
      SLAVE_LEN_WIDTH           => BUS_LEN_WIDTH,
      SLAVE_MAX_BURST           => BUS_WRITE_BURST_MAX_LEN,
      ENABLE_FIFO               => false,
      SLV_REQ_SLICE_DEPTH       => 0,
      SLV_DAT_SLICE_DEPTH       => 0,
      MST_REQ_SLICE_DEPTH       => 0,
      MST_DAT_SLICE_DEPTH       => 0
    )
    port map (
      clk                       => bus_clk,
      reset_n                   => bus_reset_n,
      slv_bus_wreq_addr         => wr_mst_wreq_addr,
      slv_bus_wreq_len          => wr_mst_wreq_len,
      slv_bus_wreq_valid        => wr_mst_wreq_valid,
      slv_bus_wreq_ready        => wr_mst_wreq_ready,
      slv_bus_wdat_data         => wr_mst_wdat_data,
      slv_bus_wdat_strobe       => wr_mst_wdat_strobe,
      slv_bus_wdat_last         => wr_mst_wdat_last,
      slv_bus_wdat_valid        => wr_mst_wdat_valid,
      slv_bus_wdat_ready        => wr_mst_wdat_ready,
      m_axi_awaddr              => m_axi_awaddr,
      m_axi_awlen               => m_axi_awlen,
      m_axi_awvalid             => m_axi_awvalid_int,
      m_axi_awready             => m_axi_awready,
      m_axi_awsize              => m_axi_awsize,
      m_axi_wdata               => m_axi_wdata,
      m_axi_wstrb               => m_axi_wstrb,
      m_axi_wlast               => m_axi_wlast,
      m_axi_wvalid              => m_axi_wvalid,
      m_axi_wready              => m_axi_wready
    );

  -- Determine the number of outstanding write requests to see if writes are
  -- pending.
  reg_proc: process (bus_clk) is
    variable outstanding  : unsigned(9 downto 0);
  begin
    if rising_edge(bus_clk) then
      write_busy <= m_axi_awvalid_int or not outstanding(9);
      if m_axi_awvalid_int = '1' and m_axi_awready = '1' then
        outstanding := outstanding + 1;
      end if;
      if m_axi_bvalid = '1' then
        outstanding := outstanding - 1;
      end if;
      if bus_reset = '1' then
        outstanding := (others => '1');
        write_busy <= '0';
      end if;
    end if;
  end process;

  m_axi_awvalid <= m_axi_awvalid_int;
  m_axi_bready <= '1';

  -----------------------------------------------------------------------------
  -- Bus arbiters
  -----------------------------------------------------------------------------
  read_arbiter_inst : entity work.BusReadArbiter
    generic map (
      BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH            => BUS_READ_INNER_DATA_WIDTH,
      NUM_SLAVE_PORTS           => 4,
      ARB_METHOD                => "RR-STICKY",
      MAX_OUTSTANDING           => 8,
      RAM_CONFIG                => "",
      SLV_REQ_SLICES            => true,
      MST_REQ_SLICE             => true,
      MST_DAT_SLICE             => true,
      SLV_DAT_SLICES            => true
    )
    port map (
      bcd_clk                   => bus_clk,
      bcd_reset                 => bus_reset,

      mst_rreq_valid            => rd_mst_rreq_valid,
      mst_rreq_ready            => rd_mst_rreq_ready,
      mst_rreq_addr             => rd_mst_rreq_addr,
      mst_rreq_len              => rd_mst_rreq_len,
      mst_rdat_valid            => rd_mst_rdat_valid,
      mst_rdat_ready            => rd_mst_rdat_ready,
      mst_rdat_data             => rd_mst_rdat_data,
      mst_rdat_last             => rd_mst_rdat_last,

      bs00_rreq_valid           => pages_text_bus_req(0).rreq_valid,
      bs00_rreq_ready           => pages_text_bus_rep(0).rreq_ready,
      bs00_rreq_addr            => pages_text_bus_req(0).rreq_addr,
      bs00_rreq_len             => pages_text_bus_req(0).rreq_len,
      bs00_rdat_valid           => pages_text_bus_rep(0).rdat_valid,
      bs00_rdat_ready           => pages_text_bus_req(0).rdat_ready,
      bs00_rdat_data            => pages_text_bus_rep(0).rdat_data,
      bs00_rdat_last            => pages_text_bus_rep(0).rdat_last,

      bs01_rreq_valid           => pages_text_bus_req(1).rreq_valid,
      bs01_rreq_ready           => pages_text_bus_rep(1).rreq_ready,
      bs01_rreq_addr            => pages_text_bus_req(1).rreq_addr,
      bs01_rreq_len             => pages_text_bus_req(1).rreq_len,
      bs01_rdat_valid           => pages_text_bus_rep(1).rdat_valid,
      bs01_rdat_ready           => pages_text_bus_req(1).rdat_ready,
      bs01_rdat_data            => pages_text_bus_rep(1).rdat_data,
      bs01_rdat_last            => pages_text_bus_rep(1).rdat_last,

      bs02_rreq_valid           => pages_text_bus_req(2).rreq_valid,
      bs02_rreq_ready           => pages_text_bus_rep(2).rreq_ready,
      bs02_rreq_addr            => pages_text_bus_req(2).rreq_addr,
      bs02_rreq_len             => pages_text_bus_req(2).rreq_len,
      bs02_rdat_valid           => pages_text_bus_rep(2).rdat_valid,
      bs02_rdat_ready           => pages_text_bus_req(2).rdat_ready,
      bs02_rdat_data            => pages_text_bus_rep(2).rdat_data,
      bs02_rdat_last            => pages_text_bus_rep(2).rdat_last,

      bs03_rreq_valid           => pages_title_bus_req.rreq_valid,
      bs03_rreq_ready           => pages_title_bus_rep.rreq_ready,
      bs03_rreq_addr            => pages_title_bus_req.rreq_addr,
      bs03_rreq_len             => pages_title_bus_req.rreq_len,
      bs03_rdat_valid           => pages_title_bus_rep.rdat_valid,
      bs03_rdat_ready           => pages_title_bus_req.rdat_ready,
      bs03_rdat_data            => pages_title_bus_rep.rdat_data,
      bs03_rdat_last            => pages_title_bus_rep.rdat_last
    );

  write_arbiter_inst : entity work.BusWriteArbiter
    generic map (
      BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH            => BUS_WRITE_INNER_DATA_WIDTH,
      NUM_SLAVE_PORTS           => 2,
      ARB_METHOD                => "RR-STICKY",
      MAX_OUTSTANDING           => 4,
      RAM_CONFIG                => "",
      SLV_REQ_SLICES            => true,
      MST_REQ_SLICE             => true,
      MST_DAT_SLICE             => true,
      SLV_DAT_SLICES            => true
    )
    port map (
      bcd_clk                   => bus_clk,
      bcd_reset                 => bus_reset,

      mst_wreq_valid            => wr_mst_wreq_valid,
      mst_wreq_ready            => wr_mst_wreq_ready,
      mst_wreq_addr             => wr_mst_wreq_addr,
      mst_wreq_len              => wr_mst_wreq_len,
      mst_wdat_valid            => wr_mst_wdat_valid,
      mst_wdat_ready            => wr_mst_wdat_ready,
      mst_wdat_data             => wr_mst_wdat_data,
      mst_wdat_strobe           => wr_mst_wdat_strobe,
      mst_wdat_last             => wr_mst_wdat_last,

      bs00_wreq_valid           => result_title_bus_req.wreq_valid,
      bs00_wreq_ready           => result_title_bus_rep.wreq_ready,
      bs00_wreq_addr            => result_title_bus_req.wreq_addr,
      bs00_wreq_len             => result_title_bus_req.wreq_len,
      bs00_wdat_valid           => result_title_bus_req.wdat_valid,
      bs00_wdat_ready           => result_title_bus_rep.wdat_ready,
      bs00_wdat_data            => result_title_bus_req.wdat_data,
      bs00_wdat_strobe          => result_title_bus_req.wdat_strobe,
      bs00_wdat_last            => result_title_bus_req.wdat_last,

      bs01_wreq_valid           => result_count_stats_bus_req.wreq_valid,
      bs01_wreq_ready           => result_count_stats_bus_rep.wreq_ready,
      bs01_wreq_addr            => result_count_stats_bus_req.wreq_addr,
      bs01_wreq_len             => result_count_stats_bus_req.wreq_len,
      bs01_wdat_valid           => result_count_stats_bus_req.wdat_valid,
      bs01_wdat_ready           => result_count_stats_bus_rep.wdat_ready,
      bs01_wdat_data            => result_count_stats_bus_req.wdat_data,
      bs01_wdat_strobe          => result_count_stats_bus_req.wdat_strobe,
      bs01_wdat_last            => result_count_stats_bus_req.wdat_last
    );

  -----------------------------------------------------------------------------
  -- Fletcher readers and decompression/match datapath
  -----------------------------------------------------------------------------
  pages_text_cmd_ctrl <= pages_text_cmd_valuesAddr & pages_text_cmd_offsetAddr;

  text_read_gen: for i in 0 to 2 generate

    -- Article text length stream. This stream is actually unused.
    signal pages_text_valid         : std_logic;
    signal pages_text_ready         : std_logic;
    signal pages_text_dvalid        : std_logic;
    signal pages_text_last          : std_logic;
    signal pages_text_length        : std_logic_vector(31 downto 0);
    signal pages_text_count         : std_logic_vector(0 downto 0);

    -- Compressed article text stream.
    signal pages_text_bytes_valid   : std_logic;
    signal pages_text_bytes_ready   : std_logic;
    signal pages_text_bytes_dvalid  : std_logic;
    signal pages_text_bytes_last    : std_logic;
    signal pages_text_bytes_data    : std_logic_vector(63 downto 0);
    signal pages_text_bytes_count   : std_logic_vector(3 downto 0);

    -- Decompressed article text stream.
    signal pages_text_chars_valid   : std_logic;
    signal pages_text_chars_ready   : std_logic;
    signal pages_text_chars_dvalid  : std_logic;
    signal pages_text_chars_last    : std_logic;
    signal pages_text_chars_data    : std_logic_vector(63 downto 0);
    signal pages_text_chars_count   : std_logic_vector(3 downto 0);

  begin

    -- Article data reader.
    pages_text_reader_inst : ArrayReader
      generic map (
        BUS_ADDR_WIDTH          => BUS_ADDR_WIDTH,
        BUS_LEN_WIDTH           => BUS_LEN_WIDTH,
        BUS_DATA_WIDTH          => BUS_READ_INNER_DATA_WIDTH,
        BUS_BURST_STEP_LEN      => BUS_READ_BURST_STEP_LEN,
        BUS_BURST_MAX_LEN       => BUS_READ_BURST_MAX_LEN,
        INDEX_WIDTH             => 32,
        CFG                     => "listprim(8;epc=8,idx_fifo_xclk_stages=2,fifo_xclk_stages=2,bus_fifo_depth=300)",
        CMD_TAG_ENABLE          => true,
        CMD_TAG_WIDTH           => 1
      )
      port map (
        bcd_clk                 => bus_clk,
        bcd_reset               => bus_reset,
        kcd_clk                 => dec_clk,
        kcd_reset               => dec_reset,

        bus_rreq_valid          => pages_text_bus_req(i).rreq_valid,
        bus_rreq_ready          => pages_text_bus_rep(i).rreq_ready,
        bus_rreq_addr           => pages_text_bus_req(i).rreq_addr,
        bus_rreq_len            => pages_text_bus_req(i).rreq_len,
        bus_rdat_valid          => pages_text_bus_rep(i).rdat_valid,
        bus_rdat_ready          => pages_text_bus_req(i).rdat_ready,
        bus_rdat_data           => pages_text_bus_rep(i).rdat_data,
        bus_rdat_last           => pages_text_bus_rep(i).rdat_last,

        cmd_valid               => pages_text_cmd_valid(i),
        cmd_ready               => pages_text_cmd_ready(i),
        cmd_firstIdx            => pages_text_cmd_idx(i*32+31 downto i*32+0),
        cmd_lastidx             => pages_text_cmd_idx(i*32+63 downto i*32+32),
        cmd_ctrl                => pages_text_cmd_ctrl,
        unl_valid               => pages_text_unl_valid(i),
        unl_ready               => pages_text_unl_ready(i),

        out_valid(1)            => pages_text_bytes_valid,
        out_valid(0)            => pages_text_valid,
        out_ready(1)            => pages_text_bytes_ready,
        out_ready(0)            => pages_text_ready,
        out_data(100 downto 97) => pages_text_bytes_count,
        out_data(96 downto 33)  => pages_text_bytes_data,
        out_data(32 downto 32)  => pages_text_count,
        out_data(31 downto 0)   => pages_text_length,
        out_dvalid(1)           => pages_text_bytes_dvalid,
        out_dvalid(0)           => pages_text_dvalid,
        out_last(1)             => pages_text_bytes_last,
        out_last(0)             => pages_text_last
      );

    -- Void the length stream; we don't need it.
    pages_text_ready <= '1';

    -- Decompress the articles.
    vhsnunzip_inst: vhsnunzip_unbuffered
      generic map (
        RAM_STYLE               => "URAM"
      )
      port map (
        clk                     => dec_clk,
        reset                   => dec_reset,

        co_valid                => pages_text_bytes_valid,
        co_ready                => pages_text_bytes_ready,
        co_data                 => pages_text_bytes_data,
        co_cnt                  => pages_text_bytes_count(2 downto 0),
        co_last                 => pages_text_bytes_last,

        de_valid                => pages_text_chars_valid,
        de_ready                => pages_text_chars_ready,
        de_dvalid               => pages_text_chars_dvalid,
        de_data                 => pages_text_chars_data,
        de_cnt                  => pages_text_chars_count,
        de_last                 => pages_text_chars_last
      );

    -- Match decompressed article text against the search pattern.
    matcher_inst: entity work.WordMatch_Matcher
      port map (
        clk                     => dec_clk,
        reset                   => dec_reset,

        mmio_cfg                => mmio_cfg, -- TODO: need false path constraint on this!

        pages_text_chars_valid  => pages_text_chars_valid,
        pages_text_chars_ready  => pages_text_chars_ready,
        pages_text_chars_dvalid => pages_text_chars_dvalid,
        pages_text_chars_last   => pages_text_chars_last,
        pages_text_chars_data   => pages_text_chars_data,
        pages_text_chars_count  => pages_text_chars_count,

        match_count_valid       => match_count_part_valid(i),
        match_count_ready       => match_count_part_ready(i),
        match_count_amount      => match_count_part_amount(i*16+15 downto i*16)
      );

  end generate;

  -- Combine the three match streams into one.
  match_count_arb_inst: entity work.StreamArb
    generic map (
      NUM_INPUTS                => 3,
      INDEX_WIDTH               => 2,
      DATA_WIDTH                => 16
    )
    port map (
      clk                       => dec_clk,
      reset                     => dec_reset,

      in_valid                  => match_count_part_valid,
      in_ready                  => match_count_part_ready,
      in_data                   => match_count_part_amount,

      out_valid                 => match_count_arb_valid,
      out_ready                 => match_count_arb_ready,
      out_data                  => match_count_arb_amount,
      out_index                 => match_count_arb_part
    );

  -- Convert the match count stream to the bus clock domain.
  match_count_xclk_inst: entity work.StreamFIFO
    generic map (
      DEPTH_LOG2                => 4,
      DATA_WIDTH                => 18,
      XCLK_STAGES               => 2,
      RAM_CONFIG                => ""
    )
    port map (
      in_clk                    => dec_clk,
      in_reset                  => dec_reset,

      in_valid                  => match_count_arb_valid,
      in_ready                  => match_count_arb_ready,
      in_data(17 downto 16)     => match_count_arb_part,
      in_data(15 downto 0)      => match_count_arb_amount,

      out_clk                   => bus_clk,
      out_reset                 => bus_reset,

      out_valid                 => match_count_xclk_valid,
      out_ready                 => match_count_xclk_ready,
      out_data(17 downto 16)    => match_count_xclk_part,
      out_data(15 downto 0)     => match_count_xclk_amount
    );

  -- Article title reader.
  pages_title_reader_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH            => BUS_READ_INNER_DATA_WIDTH,
      BUS_BURST_STEP_LEN        => BUS_READ_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN         => BUS_READ_BURST_MAX_LEN,
      INDEX_WIDTH               => 32,
      CFG                       => "listprim(8)",
      CMD_TAG_ENABLE            => true,
      CMD_TAG_WIDTH             => 1
    )
    port map (
      bcd_clk                   => bus_clk,
      bcd_reset                 => bus_reset,
      kcd_clk                   => bus_clk,
      kcd_reset                 => bus_reset,

      bus_rreq_valid            => pages_title_bus_req.rreq_valid,
      bus_rreq_ready            => pages_title_bus_rep.rreq_ready,
      bus_rreq_addr             => pages_title_bus_req.rreq_addr,
      bus_rreq_len              => pages_title_bus_req.rreq_len,
      bus_rdat_valid            => pages_title_bus_rep.rdat_valid,
      bus_rdat_ready            => pages_title_bus_req.rdat_ready,
      bus_rdat_data             => pages_title_bus_rep.rdat_data,
      bus_rdat_last             => pages_title_bus_rep.rdat_last,

      cmd_valid                 => pages_title_cmd_valid,
      cmd_ready                 => pages_title_cmd_ready,
      cmd_firstIdx              => pages_title_cmd_firstIdx,
      cmd_lastidx               => pages_title_cmd_lastidx,
      cmd_ctrl                  => pages_title_cmd_ctrl,
      unl_valid                 => pages_title_unl_valid,
      unl_ready                 => pages_title_unl_ready,

      out_valid(1)              => pages_title_chars_valid,
      out_valid(0)              => pages_title_valid,
      out_ready(1)              => pages_title_chars_ready,
      out_ready(0)              => pages_title_ready,
      out_data(41 downto 41)    => pages_title_chars_count,
      out_data(40 downto 33)    => pages_title_chars_data,
      out_data(32 downto 32)    => pages_title_count,
      out_data(31 downto 0)     => pages_title_length,
      out_dvalid(1)             => pages_title_chars_dvalid,
      out_dvalid(0)             => pages_title_dvalid,
      out_last(1)               => pages_title_chars_last,
      out_last(0)               => pages_title_last
    );

  pages_title_cmd_ctrl <= pages_title_cmd_valuesAddr & pages_title_cmd_offsetAddr;

  -----------------------------------------------------------------------------
  -- Fletcher writers
  -----------------------------------------------------------------------------
  result_title_writer_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH            => BUS_WRITE_INNER_DATA_WIDTH,
      BUS_STROBE_WIDTH          => BUS_WRITE_INNER_DATA_WIDTH/8,
      BUS_BURST_STEP_LEN        => BUS_WRITE_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN         => BUS_WRITE_BURST_MAX_LEN,
      INDEX_WIDTH               => 32,
      CFG                       => "listprim(8;last_from_length=0)",
      CMD_TAG_ENABLE            => true,
      CMD_TAG_WIDTH             => 1
    )
    port map (
      bcd_clk                   => bus_clk,
      bcd_reset                 => bus_reset,
      kcd_clk                   => bus_clk,
      kcd_reset                 => bus_reset,

      bus_wreq_valid            => result_title_bus_req.wreq_valid,
      bus_wreq_ready            => result_title_bus_rep.wreq_ready,
      bus_wreq_addr             => result_title_bus_req.wreq_addr,
      bus_wreq_len              => result_title_bus_req.wreq_len,
      bus_wdat_valid            => result_title_bus_req.wdat_valid,
      bus_wdat_ready            => result_title_bus_rep.wdat_ready,
      bus_wdat_data             => result_title_bus_req.wdat_data,
      bus_wdat_strobe           => result_title_bus_req.wdat_strobe,
      bus_wdat_last             => result_title_bus_req.wdat_last,

      cmd_valid                 => result_title_cmd_valid,
      cmd_ready                 => result_title_cmd_ready,
      cmd_firstIdx              => result_title_cmd_firstIdx,
      cmd_lastidx               => result_title_cmd_lastidx,
      cmd_ctrl                  => result_title_cmd_ctrl,
      unl_valid                 => result_title_unl_valid,
      unl_ready                 => result_title_unl_ready,

      in_valid(1)               => result_title_chars_valid,
      in_valid(0)               => result_title_valid,
      in_ready(1)               => result_title_chars_ready,
      in_ready(0)               => result_title_ready,
      in_data(41 downto 41)     => result_title_chars_count,
      in_data(40 downto 33)     => result_title_chars_data,
      in_data(32 downto 32)     => result_title_count,
      in_data(31 downto 0)      => result_title_length,
      in_dvalid(1)              => result_title_chars_dvalid,
      in_dvalid(0)              => result_title_dvalid,
      in_last(1)                => result_title_chars_last,
      in_last(0)                => result_title_last
    );

  result_title_cmd_ctrl <= result_title_cmd_valuesAddr & result_title_cmd_offsetAddr;

  result_count_stats_writer_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH            => BUS_WRITE_INNER_DATA_WIDTH,
      BUS_STROBE_WIDTH          => BUS_WRITE_INNER_DATA_WIDTH/8,
      BUS_BURST_STEP_LEN        => BUS_WRITE_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN         => BUS_WRITE_BURST_MAX_LEN,
      INDEX_WIDTH               => 32,
      CFG                       => "prim(32)",
      CMD_TAG_ENABLE            => true,
      CMD_TAG_WIDTH             => 1
    )
    port map (
      bcd_clk                   => bus_clk,
      bcd_reset                 => bus_reset,
      kcd_clk                   => bus_clk,
      kcd_reset                 => bus_reset,

      bus_wreq_valid            => result_count_stats_bus_req.wreq_valid,
      bus_wreq_ready            => result_count_stats_bus_rep.wreq_ready,
      bus_wreq_addr             => result_count_stats_bus_req.wreq_addr,
      bus_wreq_len              => result_count_stats_bus_req.wreq_len,
      bus_wdat_valid            => result_count_stats_bus_req.wdat_valid,
      bus_wdat_ready            => result_count_stats_bus_rep.wdat_ready,
      bus_wdat_data             => result_count_stats_bus_req.wdat_data,
      bus_wdat_strobe           => result_count_stats_bus_req.wdat_strobe,
      bus_wdat_last             => result_count_stats_bus_req.wdat_last,

      cmd_valid                 => result_count_stats_cmd_valid,
      cmd_ready                 => result_count_stats_cmd_ready,
      cmd_firstIdx              => result_count_stats_cmd_firstIdx,
      cmd_lastidx               => result_count_stats_cmd_lastidx,
      cmd_ctrl                  => result_count_stats_cmd_addr,
      unl_valid                 => result_count_stats_unl_valid,
      unl_ready                 => result_count_stats_unl_ready,

      in_valid(0)               => result_count_stats_valid,
      in_ready(0)               => result_count_stats_ready,
      in_data(31 downto 0)      => result_count_stats_data,
      in_dvalid(0)              => result_count_stats_dvalid,
      in_last(0)                => result_count_stats_last
    );

  -----------------------------------------------------------------------------
  -- Control logic
  -----------------------------------------------------------------------------
  cmd_gen_inst: entity work.WordMatch_CmdGen
    generic map (
      BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH
    )
    port map (
      clk                       => bus_clk,
      reset                     => bus_reset,

      mmio_cmd                  => mmio_cmd,
      mmio_start                => mmio_start,
      mmio_starting             => mmio_starting,
      mmio_done                 => mmio_done,

      pages_text_cmd_valid      => pages_text_cmd_valid,
      pages_text_cmd_ready      => pages_text_cmd_ready,
      pages_text_cmd_idx        => pages_text_cmd_idx,
      pages_text_cmd_valuesAddr => pages_text_cmd_valuesAddr,
      pages_text_cmd_offsetAddr => pages_text_cmd_offsetAddr,
      pages_text_unl_valid      => pages_text_unl_valid,
      pages_text_unl_ready      => pages_text_unl_ready,

      match_count_in_valid      => match_count_xclk_valid,
      match_count_in_ready      => match_count_xclk_ready,
      match_count_in_amount     => match_count_xclk_amount,
      match_count_in_part       => match_count_xclk_part,

      match_count_out_valid     => match_count_tagged_valid,
      match_count_out_ready     => match_count_tagged_ready,
      match_count_out_amount    => match_count_tagged_amount,
      match_count_out_index     => match_count_tagged_index,
      match_count_out_last      => match_count_tagged_last,

      result_title_cmd_valid          => result_title_cmd_valid,
      result_title_cmd_ready          => result_title_cmd_ready,
      result_title_cmd_firstIdx       => result_title_cmd_firstIdx,
      result_title_cmd_lastIdx        => result_title_cmd_lastIdx,
      result_title_cmd_valuesAddr     => result_title_cmd_valuesAddr,
      result_title_cmd_offsetAddr     => result_title_cmd_offsetAddr,
      result_title_unl_valid          => result_title_unl_valid,
      result_title_unl_ready          => result_title_unl_ready,

      result_count_stats_cmd_valid    => result_count_stats_cmd_valid,
      result_count_stats_cmd_ready    => result_count_stats_cmd_ready,
      result_count_stats_cmd_firstIdx => result_count_stats_cmd_firstIdx,
      result_count_stats_cmd_lastidx  => result_count_stats_cmd_lastidx,
      result_count_stats_cmd_addr     => result_count_stats_cmd_addr,
      result_count_stats_unl_valid    => result_count_stats_unl_valid,
      result_count_stats_unl_ready    => result_count_stats_unl_ready,

      write_busy                => write_busy
    );

  filter_inst: entity work.WordMatch_Filter
    generic map (
      BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH
    )
    port map (
      clk                       => bus_clk,
      reset                     => bus_reset,

      mmio_filt                 => mmio_filt,
      mmio_stat                 => mmio_stat,
      mmio_starting             => mmio_starting,

      match_count_valid         => match_count_tagged_valid,
      match_count_ready         => match_count_tagged_ready,
      match_count_amount        => match_count_tagged_amount,
      match_count_index         => match_count_tagged_index,
      match_count_last          => match_count_tagged_last,

      pages_title_cmd_valid     => pages_title_cmd_valid,
      pages_title_cmd_ready     => pages_title_cmd_ready,
      pages_title_cmd_firstIdx  => pages_title_cmd_firstIdx,
      pages_title_cmd_lastidx   => pages_title_cmd_lastidx,
      pages_title_cmd_valuesAddr=> pages_title_cmd_valuesAddr,
      pages_title_cmd_offsetAddr=> pages_title_cmd_offsetAddr,
      pages_title_unl_valid     => pages_title_unl_valid,
      pages_title_unl_ready     => pages_title_unl_ready,

      write_cmd_valid           => write_cmd_valid,
      write_cmd_ready           => write_cmd_ready,
      write_cmd_titlePass       => write_cmd_titlePass,
      write_cmd_titleDummy      => write_cmd_titleDummy,
      write_cmd_titleTerm       => write_cmd_titleTerm,
      write_cmd_intEnable       => write_cmd_intEnable,
      write_cmd_intData         => write_cmd_intData,
      write_cmd_last            => write_cmd_last
    );

  result_writer_inst: entity work.WordMatch_ResultWriter
    port map (
      clk                       => bus_clk,
      reset                     => bus_reset,

      write_cmd_valid           => write_cmd_valid,
      write_cmd_ready           => write_cmd_ready,
      write_cmd_titlePass       => write_cmd_titlePass,
      write_cmd_titleDummy      => write_cmd_titleDummy,
      write_cmd_titleTerm       => write_cmd_titleTerm,
      write_cmd_intEnable       => write_cmd_intEnable,
      write_cmd_intData         => write_cmd_intData,
      write_cmd_last            => write_cmd_last,

      pages_title_valid         => pages_title_valid,
      pages_title_ready         => pages_title_ready,
      pages_title_dvalid        => pages_title_dvalid,
      pages_title_last          => pages_title_last,
      pages_title_length        => pages_title_length,
      pages_title_count         => pages_title_count,
      pages_title_chars_valid   => pages_title_chars_valid,
      pages_title_chars_ready   => pages_title_chars_ready,
      pages_title_chars_dvalid  => pages_title_chars_dvalid,
      pages_title_chars_last    => pages_title_chars_last,
      pages_title_chars_data    => pages_title_chars_data,
      pages_title_chars_count   => pages_title_chars_count,

      result_title_valid        => result_title_valid,
      result_title_ready        => result_title_ready,
      result_title_dvalid       => result_title_dvalid,
      result_title_last         => result_title_last,
      result_title_length       => result_title_length,
      result_title_count        => result_title_count,
      result_title_chars_valid  => result_title_chars_valid,
      result_title_chars_ready  => result_title_chars_ready,
      result_title_chars_dvalid => result_title_chars_dvalid,
      result_title_chars_last   => result_title_chars_last,
      result_title_chars_data   => result_title_chars_data,
      result_title_chars_count  => result_title_chars_count,

      result_count_stats_valid  => result_count_stats_valid,
      result_count_stats_ready  => result_count_stats_ready,
      result_count_stats_data   => result_count_stats_data,
      result_count_stats_dvalid => result_count_stats_dvalid,
      result_count_stats_last   => result_count_stats_last
    );

end architecture;
