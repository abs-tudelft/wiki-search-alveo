library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity word_match is
  generic (
    BUS_ADDR_WIDTH : integer := 64
  );
  port (
    kcd_clk                   : in  std_logic;
    kcd_reset                 : in  std_logic;
    mmio_awvalid              : in  std_logic;
    mmio_awready              : out std_logic;
    mmio_awaddr               : in  std_logic_vector(31 downto 0);
    mmio_wvalid               : in  std_logic;
    mmio_wready               : out std_logic;
    mmio_wdata                : in  std_logic_vector(31 downto 0);
    mmio_wstrb                : in  std_logic_vector(3 downto 0);
    mmio_bvalid               : out std_logic;
    mmio_bready               : in  std_logic;
    mmio_bresp                : out std_logic_vector(1 downto 0);
    mmio_arvalid              : in  std_logic;
    mmio_arready              : out std_logic;
    mmio_araddr               : in  std_logic_vector(31 downto 0);
    mmio_rvalid               : out std_logic;
    mmio_rready               : in  std_logic;
    mmio_rdata                : out std_logic_vector(31 downto 0);
    mmio_rresp                : out std_logic_vector(1 downto 0);
    Pages_title_valid         : in  std_logic;
    Pages_title_ready         : out std_logic;
    Pages_title_dvalid        : in  std_logic;
    Pages_title_last          : in  std_logic;
    Pages_title_length        : in  std_logic_vector(31 downto 0);
    Pages_title_count         : in  std_logic_vector(0 downto 0);
    Pages_title_chars_valid   : in  std_logic;
    Pages_title_chars_ready   : out std_logic;
    Pages_title_chars_dvalid  : in  std_logic;
    Pages_title_chars_last    : in  std_logic;
    Pages_title_chars_data    : in  std_logic_vector(7 downto 0);
    Pages_title_chars_count   : in  std_logic_vector(0 downto 0);
    Pages_title_cmd_valid     : out std_logic;
    Pages_title_cmd_ready     : in  std_logic;
    Pages_title_cmd_firstIdx  : out std_logic_vector(31 downto 0);
    Pages_title_cmd_lastidx   : out std_logic_vector(31 downto 0);
    Pages_title_cmd_ctrl      : out std_logic_vector(2*bus_addr_width-1 downto 0);
    Pages_title_cmd_tag       : out std_logic_vector(0 downto 0);
    Pages_title_unl_valid     : in  std_logic;
    Pages_title_unl_ready     : out std_logic;
    Pages_title_unl_tag       : in  std_logic_vector(0 downto 0);
    Pages_text_valid          : in  std_logic;
    Pages_text_ready          : out std_logic;
    Pages_text_dvalid         : in  std_logic;
    Pages_text_last           : in  std_logic;
    Pages_text_length         : in  std_logic_vector(31 downto 0);
    Pages_text_count          : in  std_logic_vector(0 downto 0);
    Pages_text_bytes_valid    : in  std_logic;
    Pages_text_bytes_ready    : out std_logic;
    Pages_text_bytes_dvalid   : in  std_logic;
    Pages_text_bytes_last     : in  std_logic;
    Pages_text_bytes_data     : in  std_logic_vector(63 downto 0);
    Pages_text_bytes_count    : in  std_logic_vector(3 downto 0);
    Pages_text_cmd_valid      : out std_logic;
    Pages_text_cmd_ready      : in  std_logic;
    Pages_text_cmd_firstIdx   : out std_logic_vector(31 downto 0);
    Pages_text_cmd_lastidx    : out std_logic_vector(31 downto 0);
    Pages_text_cmd_ctrl       : out std_logic_vector(2*bus_addr_width-1 downto 0);
    Pages_text_cmd_tag        : out std_logic_vector(0 downto 0);
    Pages_text_unl_valid      : in  std_logic;
    Pages_text_unl_ready      : out std_logic;
    Pages_text_unl_tag        : in  std_logic_vector(0 downto 0);
    Result_title_valid        : out std_logic;
    Result_title_ready        : in  std_logic;
    Result_title_dvalid       : out std_logic;
    Result_title_last         : out std_logic;
    Result_title_length       : out std_logic_vector(31 downto 0);
    Result_title_count        : out std_logic_vector(0 downto 0);
    Result_title_chars_valid  : out std_logic;
    Result_title_chars_ready  : in  std_logic;
    Result_title_chars_dvalid : out std_logic;
    Result_title_chars_last   : out std_logic;
    Result_title_chars_data   : out std_logic_vector(7 downto 0);
    Result_title_chars_count  : out std_logic_vector(0 downto 0);
    Result_title_cmd_valid    : out std_logic;
    Result_title_cmd_ready    : in  std_logic;
    Result_title_cmd_firstIdx : out std_logic_vector(31 downto 0);
    Result_title_cmd_lastidx  : out std_logic_vector(31 downto 0);
    Result_title_cmd_ctrl     : out std_logic_vector(2*bus_addr_width-1 downto 0);
    Result_title_cmd_tag      : out std_logic_vector(0 downto 0);
    Result_title_unl_valid    : in  std_logic;
    Result_title_unl_ready    : out std_logic;
    Result_title_unl_tag      : in  std_logic_vector(0 downto 0);
    Result_count_valid        : out std_logic;
    Result_count_ready        : in  std_logic;
    Result_count_dvalid       : out std_logic;
    Result_count_last         : out std_logic;
    Result_count              : out std_logic_vector(31 downto 0);
    Result_count_cmd_valid    : out std_logic;
    Result_count_cmd_ready    : in  std_logic;
    Result_count_cmd_firstIdx : out std_logic_vector(31 downto 0);
    Result_count_cmd_lastidx  : out std_logic_vector(31 downto 0);
    Result_count_cmd_ctrl     : out std_logic_vector(bus_addr_width-1 downto 0);
    Result_count_cmd_tag      : out std_logic_vector(0 downto 0);
    Result_count_unl_valid    : in  std_logic;
    Result_count_unl_ready    : out std_logic;
    Result_count_unl_tag      : in  std_logic_vector(0 downto 0);
    Stats_stats_valid         : out std_logic;
    Stats_stats_ready         : in  std_logic;
    Stats_stats_dvalid        : out std_logic;
    Stats_stats_last          : out std_logic;
    Stats_stats               : out std_logic_vector(63 downto 0);
    Stats_stats_cmd_valid     : out std_logic;
    Stats_stats_cmd_ready     : in  std_logic;
    Stats_stats_cmd_firstIdx  : out std_logic_vector(31 downto 0);
    Stats_stats_cmd_lastidx   : out std_logic_vector(31 downto 0);
    Stats_stats_cmd_ctrl      : out std_logic_vector(bus_addr_width-1 downto 0);
    Stats_stats_cmd_tag       : out std_logic_vector(0 downto 0);
    Stats_stats_unl_valid     : in  std_logic;
    Stats_stats_unl_ready     : out std_logic;
    Stats_stats_unl_tag       : in  std_logic_vector(0 downto 0)
  );
end entity;
architecture Implementation of word_match is
begin
end architecture;
